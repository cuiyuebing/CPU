`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/05/17 19:32:19
// Design Name: 
// Module Name: left_shift
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module left_shift(
    input [31:0] A,
    input [31:0] B,
    output [31:0] C,
    output [31:0] s
    );
    //c0-c31 ??????��?????32:1 mux????????????
    wire [31:0] c0;
    wire [31:0] c1;
    wire [31:0] c2;
    wire [31:0] c3;
    wire [31:0] c4;
    wire [31:0] c5;
    wire [31:0] c6;
    wire [31:0] c7;
    wire [31:0] c8;
    wire [31:0] c9;
    wire [31:0] c10;
    wire [31:0] c11;
    wire [31:0] c12;
    wire [31:0] c13;
    wire [31:0] c14;
    wire [31:0] c15;
    wire [31:0] c16;
    wire [31:0] c17;
    wire [31:0] c18;
    wire [31:0] c19;
    wire [31:0] c20;
    wire [31:0] c21;
    wire [31:0] c22;
    wire [31:0] c23;
    wire [31:0] c24;
    wire [31:0] c25;
    wire [31:0] c26;
    wire [31:0] c27;
    wire [31:0] c28;
    wire [31:0] c29;
    wire [31:0] c30;
    wire [31:0] c31;
    
    wire low;//??
    //32????????
    parameter s0 = 32'b0;
    parameter s1 = 32'b1;
    parameter s2 = 32'b10;
    parameter s3 = 32'b11;
    parameter s4 = 32'b100;
    parameter s5 = 32'b101;
    parameter s6 = 32'b110;
    parameter s7 = 32'b111;
    parameter s8 = 32'b1000;
    parameter s9 = 32'b1001;
    parameter s10 = 32'b1010;
    parameter s11 = 32'b1011;
    parameter s12 = 32'b1100;
    parameter s13 = 32'b1101;
    parameter s14 = 32'b1110;
    parameter s15 = 32'b1111;
    parameter s16 = 32'b10000;
    parameter s17 = 32'b10001;
    parameter s18 = 32'b10010;
    parameter s19 = 32'b10011;
    parameter s20 = 32'b10100;
    parameter s21 = 32'b10101;
    parameter s22 = 32'b10110;
    parameter s23 = 32'b10111;
    parameter s24 = 32'b11000;
    parameter s25 = 32'b11001;
    parameter s26 = 32'b11010;
    parameter s27 = 32'b11011;
    parameter s28 = 32'b11100;
    parameter s29 = 32'b11101;
    parameter s30 = 32'b11110;
    parameter s31 = 32'b11111;
    //?????��??????????s
    AND_f	U0(
        .a(s0),
        .b(B),
        .co(s[0])
    );
    AND_f    U1(
        .a(s1),
        .b(B),
        .co(s[1])
    );
    AND_f    U2(
        .a(s2),
        .b(B),
        .co(s[2])
    );
    AND_f    U3(
        .a(s3),
        .b(B),
        .co(s[3])
    );
    AND_f    U4(
        .a(s4),
        .b(B),
        .co(s[4])
    );
    AND_f    U5(
        .a(s5),
        .b(B),
        .co(s[5])
    );
    AND_f    U6(
        .a(s6),
        .b(B),
        .co(s[6])
    );
    AND_f    U7(
        .a(s7),
        .b(B),
        .co(s[7])
    );
    AND_f    U8(
        .a(s8),
        .b(B),
        .co(s[8])
    );
    AND_f    U9(
        .a(s9),
        .b(B),
        .co(s[9])
    );
    AND_f    U10(
        .a(s10),
        .b(B),
        .co(s[10])
    );
    AND_f    U11(
        .a(s11),
        .b(B),
        .co(s[11])
    );
    AND_f    U12(
        .a(s12),
        .b(B),
        .co(s[12])
    );
    AND_f    U13(
        .a(s13),
        .b(B),
        .co(s[13])
    );
    AND_f    U14(
        .a(s14),
        .b(B),
        .co(s[14])
    );
    AND_f    U15(
        .a(s15),
        .b(B),
        .co(s[15])
    );
    AND_f    U16(
        .a(s16),
        .b(B),
        .co(s[16])
    );
    AND_f    U17(
        .a(s17),
        .b(B),
        .co(s[17])
    );
    AND_f    U18(
        .a(s18),
        .b(B),
        .co(s[18])
    );
    AND_f    U19(
        .a(s19),
        .b(B),
        .co(s[19])
    );
    AND_f    U20(
        .a(s20),
        .b(B),
        .co(s[20])
    );
    AND_f    U21(
        .a(s21),
        .b(B),
        .co(s[21])
    );
    AND_f    U22(
        .a(s22),
        .b(B),
        .co(s[22])
    );
    AND_f    U23(
        .a(s23),
        .b(B),
        .co(s[23])
    );
    AND_f    U24(
        .a(s24),
        .b(B),
        .co(s[24])
    );
    AND_f    U25(
        .a(s25),
        .b(B),
        .co(s[25])
    );
    AND_f    U26(
        .a(s26),
        .b(B),
        .co(s[26])
    );
    AND_f    U27(
        .a(s27),
        .b(B),
        .co(s[27])
    );
    AND_f    U28(
        .a(s28),
        .b(B),
        .co(s[28])
    );
    AND_f    U29(
        .a(s29),
        .b(B),
        .co(s[29])
    );
    AND_f    U30(
        .a(s30),
        .b(B),
        .co(s[30])
    );
    AND_f    U31(
        .a(s31),
        .b(B),
        .co(s[31])
    );
    //????32??mux ????????????????
    genvar i;
    generate  
        //32:1mux *32
        for (i=0;i<32;i=i+1)
        begin
            and (c31[i], s[i], A[31 - i]);
        end
        for (i=0;i<31;i=i+1)
        begin
            and (c30[i], s[i], A[30 - i]);
        end
        for (i=0;i<30;i=i+1)
        begin
            and (c29[i], s[i], A[29 - i]);
        end
        for (i=0;i<29;i=i+1)
        begin
            and (c28[i], s[i], A[28 - i]);
        end
        for (i=0;i<28;i=i+1)
        begin
            and (c27[i], s[i], A[27 - i]);
        end
        for (i=0;i<27;i=i+1)
        begin
            and (c26[i], s[i], A[26 - i]);
        end
        for (i=0;i<26;i=i+1)
        begin
            and (c25[i], s[i], A[25 - i]);
        end
        for (i=0;i<25;i=i+1)
        begin
            and (c24[i], s[i], A[24 - i]);
        end
        for (i=0;i<24;i=i+1)
        begin
            and (c23[i], s[i], A[23 - i]);
        end
        for (i=0;i<23;i=i+1)
        begin
            and (c22[i], s[i], A[22 - i]);
        end
        for (i=0;i<22;i=i+1)
        begin
            and (c21[i], s[i], A[21 - i]);
        end
        for (i=0;i<21;i=i+1)
        begin
            and (c20[i], s[i], A[20 - i]);
        end
        for (i=0;i<20;i=i+1)
        begin
            and (c19[i], s[i], A[19 - i]);
        end
        for (i=0;i<19;i=i+1)
        begin
            and (c18[i], s[i], A[18 - i]);
        end
        for (i=0;i<18;i=i+1)
        begin
            and (c17[i], s[i], A[17 - i]);
        end
        for (i=0;i<17;i=i+1)
        begin
            and (c16[i], s[i], A[16 - i]);
        end
        for (i=0;i<16;i=i+1)
        begin
            and (c15[i], s[i], A[15 - i]);
        end
        for (i=0;i<15;i=i+1)
        begin
            and (c14[i], s[i], A[14 - i]);
        end
        for (i=0;i<14;i=i+1)
        begin
            and (c13[i], s[i], A[13 - i]);
        end
        for (i=0;i<13;i=i+1)
        begin
            and (c12[i], s[i], A[12 - i]);
        end
        for (i=0;i<12;i=i+1)
        begin
            and (c11[i], s[i], A[11 - i]);
        end
        for (i=0;i<11;i=i+1)
        begin
            and (c10[i], s[i], A[10 - i]);
        end
        for (i=0;i<10;i=i+1)
        begin
            and (c9[i], s[i], A[9 - i]);
        end
        for (i=0;i<9;i=i+1)
        begin
            and (c8[i], s[i], A[8 - i]);
        end
        for (i=0;i<8;i=i+1)
        begin
            and (c7[i], s[i], A[7 - i]);
        end
        for (i=0;i<7;i=i+1)
        begin
            and (c6[i], s[i], A[6 - i]);
        end
        for (i=0;i<6;i=i+1)
        begin
            and (c5[i], s[i], A[5 - i]);
        end
        for (i=0;i<5;i=i+1)
        begin
            and (c4[i], s[i], A[4 - i]);
        end
        for (i=0;i<4;i=i+1)
        begin
            and (c3[i], s[i], A[3 - i]);
        end
        for (i=0;i<3;i=i+1)
        begin
            and (c2[i], s[i], A[2 - i]);
        end
        for (i=0;i<2;i=i+1)
        begin
            and (c1[i], s[i], A[1 - i]);
        end
        for (i=0;i<1;i=i+1)
        begin
            and (c0[i], s[i], A[0 - i]);
        end 
    endgenerate
    
    assign low=0;//??
    //????????����??
    or (C[0],c0[0],low);
    or (C[1],c1[0],c1[1]);
    or (C[2],c2[0],c2[1],c2[2]);
    or (C[3],c3[0],c3[1],c3[2],c3[3]);
    or (C[4],c4[0],c4[1],c4[2],c4[3],c4[4]);
    or (C[5],c5[0],c5[1],c5[2],c5[3],c5[4],c5[5]);
    or (C[6],c6[0],c6[1],c6[2],c6[3],c6[4],c6[5],c6[6]);
    or (C[7],c7[0],c7[1],c7[2],c7[3],c7[4],c7[5],c7[6],c7[7]);
    or (C[8],c8[0],c8[1],c8[2],c8[3],c8[4],c8[5],c8[6],c8[7],c8[8]);
    or (C[9],c9[0],c9[1],c9[2],c9[3],c9[4],c9[5],c9[6],c9[7],c9[8],c9[9]);
    or (C[10],c10[0],c10[1],c10[2],c10[3],c10[4],c10[5],c10[6],c10[7],c10[8],c10[9],c10[10]);
    or (C[11],c11[0],c11[1],c11[2],c11[3],c11[4],c11[5],c11[6],c11[7],c11[8],c11[9],c11[10],c11[11]);
    or (C[12],c12[0],c12[1],c12[2],c12[3],c12[4],c12[5],c12[6],c12[7],c12[8],c12[9],c12[10],c12[11],c12[12]);
    or (C[13],c13[0],c13[1],c13[2],c13[3],c13[4],c13[5],c13[6],c13[7],c13[8],c13[9],c13[10],c13[11],c13[12],c13[13]);
    or (C[14],c14[0],c14[1],c14[2],c14[3],c14[4],c14[5],c14[6],c14[7],c14[8],c14[9],c14[10],c14[11],c14[12],c14[13],c14[14]);
    or (C[15],c15[0],c15[1],c15[2],c15[3],c15[4],c15[5],c15[6],c15[7],c15[8],c15[9],c15[10],c15[11],c15[12],c15[13],c15[14],c15[15]);
    or (C[16],c16[0],c16[1],c16[2],c16[3],c16[4],c16[5],c16[6],c16[7],c16[8],c16[9],c16[10],c16[11],c16[12],c16[13],c16[14],c16[15],c16[16]);
    or (C[17],c17[0],c17[1],c17[2],c17[3],c17[4],c17[5],c17[6],c17[7],c17[8],c17[9],c17[10],c17[11],c17[12],c17[13],c17[14],c17[15],c17[16],c17[17]);
    or (C[18],c18[0],c18[1],c18[2],c18[3],c18[4],c18[5],c18[6],c18[7],c18[8],c18[9],c18[10],c18[11],c18[12],c18[13],c18[14],c18[15],c18[16],c18[17],c18[18]);
    or (C[19],c19[0],c19[1],c19[2],c19[3],c19[4],c19[5],c19[6],c19[7],c19[8],c19[9],c19[10],c19[11],c19[12],c19[13],c19[14],c19[15],c19[16],c19[17],c19[18],c19[19]);
    or (C[20],c20[0],c20[1],c20[2],c20[3],c20[4],c20[5],c20[6],c20[7],c20[8],c20[9],c20[10],c20[11],c20[12],c20[13],c20[14],c20[15],c20[16],c20[17],c20[18],c20[19],c20[20]);
    or (C[21],c21[0],c21[1],c21[2],c21[3],c21[4],c21[5],c21[6],c21[7],c21[8],c21[9],c21[10],c21[11],c21[12],c21[13],c21[14],c21[15],c21[16],c21[17],c21[18],c21[19],c21[20],c21[21]);
    or (C[22],c22[0],c22[1],c22[2],c22[3],c22[4],c22[5],c22[6],c22[7],c22[8],c22[9],c22[10],c22[11],c22[12],c22[13],c22[14],c22[15],c22[16],c22[17],c22[18],c22[19],c22[20],c22[21],c22[22]);
    or (C[23],c23[0],c23[1],c23[2],c23[3],c23[4],c23[5],c23[6],c23[7],c23[8],c23[9],c23[10],c23[11],c23[12],c23[13],c23[14],c23[15],c23[16],c23[17],c23[18],c23[19],c23[20],c23[21],c23[22],c23[23]);
    or (C[24],c24[0],c24[1],c24[2],c24[3],c24[4],c24[5],c24[6],c24[7],c24[8],c24[9],c24[10],c24[11],c24[12],c24[13],c24[14],c24[15],c24[16],c24[17],c24[18],c24[19],c24[20],c24[21],c24[22],c24[23],c24[24]);
    or (C[25],c25[0],c25[1],c25[2],c25[3],c25[4],c25[5],c25[6],c25[7],c25[8],c25[9],c25[10],c25[11],c25[12],c25[13],c25[14],c25[15],c25[16],c25[17],c25[18],c25[19],c25[20],c25[21],c25[22],c25[23],c25[24],c25[25]);
    or (C[26],c26[0],c26[1],c26[2],c26[3],c26[4],c26[5],c26[6],c26[7],c26[8],c26[9],c26[10],c26[11],c26[12],c26[13],c26[14],c26[15],c26[16],c26[17],c26[18],c26[19],c26[20],c26[21],c26[22],c26[23],c26[24],c26[25],c26[26]);
    or (C[27],c27[0],c27[1],c27[2],c27[3],c27[4],c27[5],c27[6],c27[7],c27[8],c27[9],c27[10],c27[11],c27[12],c27[13],c27[14],c27[15],c27[16],c27[17],c27[18],c27[19],c27[20],c27[21],c27[22],c27[23],c27[24],c27[25],c27[26],c27[27]);
    or (C[28],c28[0],c28[1],c28[2],c28[3],c28[4],c28[5],c28[6],c28[7],c28[8],c28[9],c28[10],c28[11],c28[12],c28[13],c28[14],c28[15],c28[16],c28[17],c28[18],c28[19],c28[20],c28[21],c28[22],c28[23],c28[24],c28[25],c28[26],c28[27],c28[28]);
    or (C[29],c29[0],c29[1],c29[2],c29[3],c29[4],c29[5],c29[6],c29[7],c29[8],c29[9],c29[10],c29[11],c29[12],c29[13],c29[14],c29[15],c29[16],c29[17],c29[18],c29[19],c29[20],c29[21],c29[22],c29[23],c29[24],c29[25],c29[26],c29[27],c29[28],c29[29]);
    or (C[30],c30[0],c30[1],c30[2],c30[3],c30[4],c30[5],c30[6],c30[7],c30[8],c30[9],c30[10],c30[11],c30[12],c30[13],c30[14],c30[15],c30[16],c30[17],c30[18],c30[19],c30[20],c30[21],c30[22],c30[23],c30[24],c30[25],c30[26],c30[27],c30[28],c30[29],c30[30]);
    or (C[31],c31[0],c31[1],c31[2],c31[3],c31[4],c31[5],c31[6],c31[7],c31[8],c31[9],c31[10],c31[11],c31[12],c31[13],c31[14],c31[15],c31[16],c31[17],c31[18],c31[19],c31[20],c31[21],c31[22],c31[23],c31[24],c31[25],c31[26],c31[27],c31[28],c31[29],c31[30],c31[31]);
    
endmodule
